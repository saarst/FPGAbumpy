// (c) Technion IIT, Department of Electrical Engineering 2018 
// Written By David Bar-On  June 2018 
// detect a key and generate three ouptputs for this key 


module key_risingEdge 	
 ( 
   input	 logic     clk,
	input	 logic     resetN,
	input  logic     key,
	  
   output logic  keyRisingEdgePulse	//  valid for one clock after presing the key 
 	 
  ) ;
 
 	
	logic keyIsPressed_d,keyIsPressed ; //  _d == delay of one clock 

   assign keyRisingEdgePulse = ( keyIsPressed_d == 1'b0 ) && ( keyIsPressed == 1'b1 ) ; // detects a rising edge (change) in the input
 
  
	always_ff @(posedge clk or negedge resetN)
		begin
			if (!resetN ) begin 
				keyIsPressed_d <= 0  ; 
				keyIsPressed  <= 0 ; 
	 
			end
			
			else begin
			keyIsPressed_d  <= keyIsPressed; // generate a delay of one clock
			
			if (!key)    keyIsPressed <= 1'b1 ; 
			else 			 keyIsPressed <= 1'b0 ; 
			end  
			
			
	end // always_ff 
	

endmodule


